module viewport

import gg
import ui
import ui.component { gg_canvaslayout }
import artemkakun.trnsfrm2d

const viewport_z_index = 1

// ViewportApp is a `gg` app that represents a viewport for sprite rendering and polygon shape editing.
pub struct ViewportApp {
mut:
	gg             &gg.Context
	bounds         gg.Rect
	work_sprite    ?gg.Image
	polygon_points []trnsfrm2d.Position
}

fn (mut app ViewportApp) on_init() {
	app.set_bounds(app.bounds)
}

fn (mut app ViewportApp) on_draw() {
	app.gg.draw_rect(app.bounds.x, app.bounds.y, app.bounds.width, app.bounds.height,
		gg.Color{
		r: 211
		g: 211
		b: 211
	})

	if app.work_sprite != none {
		sprite_to_draw := app.work_sprite or { return }

		scale := 20
		sprite_width := sprite_to_draw.width * scale
		sprite_height := sprite_to_draw.height * scale

		viewport_center_x := app.bounds.x + app.bounds.width / 2
		viewport_center_y := app.bounds.y + app.bounds.height / 2

		sprite_x := viewport_center_x - sprite_width / 2
		sprite_y := viewport_center_y - sprite_height / 2

		app.gg.draw_image_by_id(sprite_x, sprite_y, sprite_width, sprite_height, sprite_to_draw.id)
	}

	for point_index, point_position in app.polygon_points {
		if point_index == app.polygon_points.len - 1 {
			app.gg.draw_line_with_config(f32(point_position.x), f32(point_position.y),
				f32(app.polygon_points[0].x), f32(app.polygon_points[0].y), gg.PenConfig{
				color: gg.Color{
					r: 0
					g: 139
					b: 139
				}
				thickness: 2
			})
		} else {
			app.gg.draw_line_with_config(f32(point_position.x), f32(point_position.y),
				f32(app.polygon_points[point_index + 1].x), f32(app.polygon_points[point_index + 1].y),
				gg.PenConfig{
				color: gg.Color{
					r: 0
					g: 139
					b: 139
				}
				thickness: 2
			})
		}
	}

	for point_position in app.polygon_points {
		app.gg.draw_circle_filled(f32(point_position.x), f32(point_position.y), 5, gg.Color{
			r: 0
			g: 255
			b: 255
		})
	}
}

fn (mut app ViewportApp) on_delegate(event &gg.Event) {
	if event.typ == .mouse_down {
		app.polygon_points << trnsfrm2d.Position{
			x: event.mouse_x
			y: event.mouse_y
		}
	}
}

fn (mut app ViewportApp) set_bounds(bb gg.Rect) {
	app.bounds = bb
}

fn (mut app ViewportApp) run() {
	app.gg.run()
}

// create_viewport_widget creates viewport canvas widget for sprite rendering and polygon shape editing.
pub fn create_viewport_widget(viewport_app &ViewportApp) &ui.CanvasLayout {
	return gg_canvaslayout(
		app: viewport_app
		z_index: viewport.viewport_z_index
	)
}

// create_viewport_app creates a new `ViewportApp` instance and returns a reference to it.
pub fn create_viewport_app() &ViewportApp {
	mut viewport_app := &ViewportApp{
		gg: unsafe { nil }
	}

	viewport_app.gg = gg.new_context(
		user_data: viewport_app
		ui_mode: true
	)

	return viewport_app
}

// open_work_sprite opens a sprite from the provided path for editing in the viewport.
pub fn (mut app ViewportApp) open_work_sprite(path_to_sprite string) ! {
	app.work_sprite = app.gg.create_image(path_to_sprite)!
}
