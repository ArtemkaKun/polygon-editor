module main

import artemkakun.ui
import app

fn main() {
	ui.run(app.create_app())
}
