module main

import app
import ui

fn main() {
	ui.run(app.create_app())
}
